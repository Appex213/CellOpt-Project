VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO DLY_CAP_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY_CAP_X1 0 0 ;
  SIZE 1 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.045 -0.15 1.045 0.15 ;
        RECT 0.775 -0.15 0.945 0.32 ;
        RECT 0.055 -0.15 0.225 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.85 0.825 0.95 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.045 1.65 1.045 1.95 ;
        RECT 0.81 1.24 0.91 1.95 ;
        RECT 0.09 1.24 0.19 1.95 ;
    END
  END VDD
  PROPERTY CatenaDesignType "deviceLevel" ;
END DLY_CAP_X1

MACRO DLY_CAP_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY_CAP_X2 0 0 ;
  SIZE 1 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.045 -0.15 1.045 0.15 ;
        RECT 0.775 -0.15 0.945 0.32 ;
        RECT 0.055 -0.15 0.225 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.85 0.825 0.95 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.045 1.65 1.045 1.95 ;
        RECT 0.81 1.24 0.91 1.95 ;
        RECT 0.09 1.24 0.19 1.95 ;
    END
  END VDD
  PROPERTY CatenaDesignType "deviceLevel" ;
END DLY_CAP_X2

MACRO DLY_CAP_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY_CAP_X4 0 0 ;
  SIZE 1 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.045 -0.15 1.045 0.15 ;
        RECT 0.775 -0.15 0.945 0.32 ;
        RECT 0.055 -0.15 0.225 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.85 0.825 0.95 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.045 1.65 1.045 1.95 ;
        RECT 0.81 1.24 0.91 1.95 ;
        RECT 0.09 1.24 0.19 1.95 ;
    END
  END VDD
  PROPERTY CatenaDesignType "deviceLevel" ;
END DLY_CAP_X4

MACRO DLY_CAP_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY_CAP_X8 0 0 ;
  SIZE 1 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.045 -0.15 1.045 0.15 ;
        RECT 0.775 -0.15 0.945 0.32 ;
        RECT 0.055 -0.15 0.225 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.85 0.825 0.95 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.045 1.65 1.045 1.95 ;
        RECT 0.81 1.24 0.91 1.95 ;
        RECT 0.09 1.24 0.19 1.95 ;
    END
  END VDD
  PROPERTY CatenaDesignType "deviceLevel" ;
END DLY_CAP_X8

END LIBRARY
